-- Multiple high frequency clocks generated using Spartan 6 FPGA
--
-- Author : Jungho Park
-- Date : November 2016
--
-- Board : Xilinx X-SP6-X9 mini board (as shown in the picture)
-- Resources for the mini board
-- http://bravelearn.com/tag/x-sp6-x9/
-- https://artofcircuits.com/product/spartan-6-fpga-development-board-xc6slx9-tqg144
--
-- Using FPGA, multiple high frequency clock signals can be generated.
-- Xilinx Spartan-6 XC6SLX9-TQG144 speed grade 2 is used for this purpose.
-- Since FPGA does not have a fixed hardware structure, it can provide
-- very wide parallel processing. In this example, I simultaneously generated
-- 8 different clock frequencies but it can be easily expanded to 100 different
-- clock frequencies. FPGA is also beneficial to clock generation because 
-- FPGA instructions are hardware operations executed at fixed cycles. 
-- Thus, clock jitter can be minimized.
-- 
-- Spartan-6 core has a PLL which can generate a very high frequency clocks 
-- (825 Mhz) as a source clock using a primary clock (50MHz).
-- The following 6 clocks are generated using the Digital Clocking Wizard.
-- The xc6slx9 is stable up to 275MHz. These clocks are used to generate
-- additional clocks using counters.
-- In this example, Clk_Out(6)(13.75MHz) is generated by dividing CLK_OUT1
-- (275MHz) by 20. Clk_Out(7)(14.7321 MHz) is generated by dividing CLK_OUT5
-- (117.857 MHz) by 8. Clk_Out(7) (14.7321MHz) can be used for a clock source
-- (14.7456 MHz) for RS232C. 
------------------------------------------------------------------------------
-- "Output    Output      Phase     Duty      Pk-to-Pk        Phase"
-- "Clock    Freq (MHz) (degrees) Cycle (%) Jitter (ps)  Error (ps)"
------------------------------------------------------------------------------
-- CLK_OUT1___275.000______0.000______50.0______203.096____221.936
-- CLK_OUT2___206.250______0.000______50.0______212.097____221.936
-- CLK_OUT3___165.000______0.000______50.0______219.401____221.936
-- CLK_OUT4___137.500______0.000______50.0______226.445____221.936
-- CLK_OUT5___117.857______0.000______50.0______234.235____221.936
-- CLK_OUT6___103.125______0.000______50.0______241.539____221.936
--
------------------------------------------------------------------------------
-- "Input Clock   Freq (MHz)    Input Jitter (UI)"
------------------------------------------------------------------------------
-- __primary__________50.000____________0.010
-- 
-- If you install another oscillator on the board (P127), you can
-- generate a different set of clocks. 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
Library UNISIM;
use UNISIM.vcomponents.all;

entity clock_pll_275MHz is

port(clk      :in std_logic;  --CLK 50M INPUT PIN 126
     --  You can also have multiple clock outputs
     clk_out :out std_logic_vector(7 downto 0); -- clock output 0 (275 MHz) Pin 115
     -- Clock output 1 (206.25 MHz) Pin 116
     -- Clock output 2 (165 MHz) Pin 117
     -- Clock output 3 (137.5 MHz) Pin 118
     -- Clock output 4 (117.857 MHz) Pin 119
     -- Clock output 5 (103.125 MHz) Pin 120
     -- Clock output 6 (13.75 MHz) Pin 121
     -- Clock output 7 (14.732 MHz) Pin 123
     miao_out :out std_logic);  -- LED OUTPUT  led display PIN 45
	  
end clock_pll_275MHz;

architecture Behavioral of clock_pll_275MHz is
  -- Number of PLL clock outputs
  constant NUM_CLK : integer := 6;
  
  -- declaration of internal clocks
  signal clk_int : std_logic_vector(5 downto 0);
  
  -- inverted clock signals
  signal clk_int_inv : std_logic_vector(5 downto 0);
  -- ODDR2 port definitions
  signal Q : std_logic;
  signal C0 : std_logic;
  signal C1 : std_logic;
  signal CE : std_logic;
  signal D0 : std_logic;
  signal D1 : std_logic;
  signal R : std_logic;
  signal S : std_logic;

-- The definition of the PLL clock generated using the Clock Wizard (pll_clock.xco)
component pll_clock
port
 (-- Clock in ports
  CLK_IN1           : in     std_logic;
  -- Clock out ports
  CLK_OUT1          : out    std_logic;
  CLK_OUT2          : out    std_logic;
  CLK_OUT3          : out    std_logic;
  CLK_OUT4          : out    std_logic;
  CLK_OUT5          : out    std_logic;
  CLK_OUT6          : out    std_logic
 );
end component;

begin
  -- Define the inverted clocks here.
  clk_int_inv <= not(clk_int);
  
  -- ODDR2: Output Double Data Rate Output Register with Set, Reset
  -- and Clock Enable.
  -- Spartan-6
  -- Xilinx HDL Libraries Guide, version 14.7
  -- internal clock signals cannot directly drive a port.
  -- So, the internal clock signal should be sent to ODDR2
  -- and ODDR2 drives the output port.
  -- ODDR2 ports for output
  gen_outclk_oddr: 
  for index in 0 to (NUM_CLK - 1) generate 
    begin
      clkout : ODDR2
      generic map(
        DDR_ALIGNMENT => "None", -- Sets output alignment to "NONE", "C0", "C1"
        INIT => '0', -- Sets initial state of the Q output to '0' or '1'
        SRTYPE => "SYNC") -- Specifies "SYNC" or "ASYNC" set/reset
      port map (
        Q => clk_out(index), -- 1-bit output data
        C0 => clk_int(index), -- 1-bit clock input
        C1 => clk_int_inv(index), -- 1-bit clock input
        CE => '1', -- 1-bit clock enable input
        D0 => '1', -- 1-bit data input (associated with C0)
        D1 => '0', -- 1-bit data input (associated with C1)
        R => '0', -- 1-bit reset input
        S => '0' -- 1-bit set input
      );
    end generate;
  
  -- The PLL clock generated using the Clock Wizard (pll_clock.xco)
  my_new_clock : pll_clock
  port map
  (-- Clock in ports
    CLK_IN1 => CLK,
    -- map clock out ports to clock internal (clk_int)
    CLK_OUT1 => clk_int(0),
    CLK_OUT2 => clk_int(1),
	 CLK_OUT3 => clk_int(2),
    CLK_OUT4 => clk_int(3),
    CLK_OUT5 => clk_int(4),
    CLK_OUT6 => clk_int(5)
  );
  
  -- define tasks to divide the clock and produce the output clock
  -- process using clk_int(0) (275 MHz)
  process(clk_int(0))
    -- defintion for counters
    variable cnt1:integer range 0 to 68749999; --frequency division by 137 500 000 (0.5 sec)
    variable cnt2:integer range 0 to 9;  --frequency division by 20
    -- flipflops
    variable ff1:std_logic; 
    variable ff2:std_logic; 
    begin
      if clk_int(0)'event and clk_int(0)='1' then
	     -- divide the clock by 137 500 000 (0.5 sec)
        if cnt1<68749999 then
          cnt1:=cnt1+1;
        else
          cnt1:=0;
          ff1:=not ff1; -- flip the flipflop
        end if;
	     -- divide the clock by 20
        if cnt2<9 then
          cnt2:=cnt2+1;
        else
          cnt2:=0;
          ff2:=not ff2; -- flip the flipflop
        end if;
      end if;
		-- blinking LED (D7) twice per second
      miao_out <= not ff1; -- output for LED
      clk_out(6) <= not ff2; -- output for Custom7 clock
    end process;

  -- process using clk_int(4) (117.857 MHz)
  process(clk_int(4))
    variable cnt1:integer range 0 to 3; -- divide the clock by 8
    variable ff1:std_logic; 
    begin
      if clk_int(4)'event and clk_int(4)='1' then
	     -- divide the clock by 8
        if cnt1<3 then
          cnt1:=cnt1+1;
        else
          cnt1:=0;
          ff1:=not ff1; -- flip the flipflop
        end if;
      end if;
	   clk_out(7) <= not ff1; -- output for Custom8 clock
    end process;
	 
end Behavioral;
